//------------------------------------------------------------------------------
// Watchdog Timer (WDT) with APB Interface
//
// Detailed Description:
// - Provides APB-accessible registers for control, timeout configuration,
//   status, feeding, and interrupt management.
// - Implements a configurable timeout counter with optional windowed mode.
// - Generates a pre-timeout interrupt and a reset signal upon timeout.
// - Supports debug mode pause and a basic clock gating mechanism for low-power operation.
//
// Abbreviations:
//  WDT      - Watchdog Timer
//  APB      - Advanced Peripheral Bus
//  PCLK     - Peripheral Clock
//  PSEL     - Peripheral Select
//  PENABLE  - Peripheral Enable
//  PWRITE   - Peripheral Write (0 = read, 1 = write)
//  PADDR    - Peripheral Address
//  PWDATA   - Peripheral Write Data
//  PRDATA   - Peripheral Read Data
//  PREADY   - Peripheral Ready
//  PSLVERR  - Peripheral Slave Error
//------------------------------------------------------------------------------

module wdt_apb (
    // APB Interface signals
    input  logic         pclk,      // APB clock
    input  logic         presetn,   // Active low reset
    input  logic         psel,      // APB peripheral select
    input  logic         penable,   // APB enable
    input  logic         pwrite,    // APB write (1) / read (0) indicator
    input  logic [7:0]   paddr,     // APB address (word-aligned)
    input  logic [31:0]  pwdata,    // APB write data
    output logic [31:0]  prdata,    // APB read data
    output logic         pready,    // APB ready signal
    output logic         pslverr,   // APB slave error signal

    // Watchdog outputs
    output logic         wdt_reset, // System reset signal generated by WDT
    output logic         wdt_int,   // Interrupt signal generated by WDT

    // External debug mode signal (active high) to pause watchdog counter
    input  logic         debug_mode
);

  //-------------------------------------------------------------------------
  // Register Address Map (word offsets)
  //-------------------------------------------------------------------------
  localparam ADDR_WDT_CTRL     = 8'h00;
  localparam ADDR_WDT_TIMEOUT  = 8'h04;
  localparam ADDR_WDT_STATUS   = 8'h08;
  localparam ADDR_WDT_FEED     = 8'h0C;
  localparam ADDR_WDT_INT_EN   = 8'h10;
  localparam ADDR_WDT_INT_STAT = 8'h14;

  //-------------------------------------------------------------------------
  // WDT_CTRL bit definitions (within 32-bit register)
  //-------------------------------------------------------------------------
  localparam CTRL_ENABLE      = 0;  // Bit 0: WDT Enable (1 = enabled)
  localparam CTRL_WINDOW_EN   = 1;  // Bit 1: Enable Windowed Mode (1 = window mode active)
  localparam CTRL_DEBUG_PAUSE = 2;  // Bit 2: Pause in Debug Mode (1 = pause)
  localparam CTRL_RESET_TYPE  = 3;  // Bit 3: Reset Type (0 = soft, 1 = hard)
  localparam CTRL_CLK_GATE    = 4;  // Bit 4: Clock Gating Enable (1 = enabled)

  //-------------------------------------------------------------------------
  // Internal registers for APB registers
  //-------------------------------------------------------------------------
  logic [31:0] reg_wdt_ctrl;
  logic [31:0] reg_wdt_timeout;
  logic [31:0] reg_wdt_status;
  logic [31:0] reg_wdt_int_en;
  logic [31:0] reg_wdt_int_stat;

  // Internal counter register (32-bit counter)
  logic [31:0] counter;

  // Parameter: Interrupt margin (number of cycles before timeout when interrupt is generated)
  localparam logic [31:0] INT_MARGIN = 32'd10;

  //-------------------------------------------------------------------------
  // Feed event: Occurs when a write to the WDT_FEED register happens AND,
  // if windowed mode is enabled, the current counter is within the valid window.
  // In non-windowed mode the feed is always accepted.
  //-------------------------------------------------------------------------
  wire feed_event;
  wire window_valid;
  assign window_valid = (reg_wdt_ctrl[CTRL_WINDOW_EN]) ? (counter >= (reg_wdt_timeout >> 1)) : 1'b1;
  assign feed_event  = psel & penable & pwrite & (paddr == ADDR_WDT_FEED) & window_valid;
  
  //-------------------------------------------------------------------------
  // Clock Gating for the Watchdog Counter
  // A simple latch-based clock gating scheme is implemented.
  // Note: In a real design, use a dedicated clock gating cell.
  //-------------------------------------------------------------------------
  logic         gate_en;
  logic         Latch_Out;
  logic         gated_clk;
  
  assign gate_en = reg_wdt_ctrl[CTRL_CLK_GATE]; // Enable gating if bit is set
  
  // A level-sensitive latch: capture the gating enable signal when pclk is low.
  always @(pclk or gate_en) begin
    if (!pclk) begin
      Latch_Out <= gate_en;
    end
  end
  
  // The gated clock is produced by ANDing the APB clock with the latch output.
  assign gated_clk = pclk && Latch_Out;
  
  // Select the clock for the counter: use gated clock when clock gating is enabled,
  // otherwise use the full APB clock.
  logic clk_counter;
  assign clk_counter = (reg_wdt_ctrl[CTRL_CLK_GATE]) ? gated_clk : pclk;

  //-------------------------------------------------------------------------
  // APB Interface: Write operations
  //-------------------------------------------------------------------------
  always_ff @(posedge pclk or negedge presetn) begin
    if (!presetn) begin
      reg_wdt_ctrl     <= 32'd0;
      reg_wdt_timeout  <= 32'd1000; // Default timeout (can be adjusted)
      reg_wdt_int_en   <= 32'd0;
      reg_wdt_int_stat <= 32'd0;
    end else begin
      if (psel & penable & pwrite) begin
        case (paddr)
          ADDR_WDT_CTRL: begin
            // Writing to WDT_CTRL updates control features including enable, window mode,
            // debug pause, reset type, and clock gating.
            reg_wdt_ctrl <= pwdata;
          end
          ADDR_WDT_TIMEOUT: begin
            // Update timeout value
            reg_wdt_timeout <= pwdata;
          end
          // Writing to the feed register resets the counter (if within a valid window)
          ADDR_WDT_FEED: begin
            // Clear any pending interrupt flag on feed
            reg_wdt_int_stat[0] <= 1'b0;
          end
          ADDR_WDT_INT_EN: begin
            // Update the interrupt enable mask
            reg_wdt_int_en <= pwdata;
          end
          // W1C: Writing '1' clears the corresponding interrupt status bit.
          ADDR_WDT_INT_STAT: begin
            reg_wdt_int_stat[0] <= reg_wdt_int_stat[0] & ~pwdata[0];
          end
          default: ; // For undefined addresses, no operation (PSLVERR will be flagged in read)
        endcase
      end
    end
  end

  //-------------------------------------------------------------------------
  // APB Interface: Read operations
  //-------------------------------------------------------------------------
  always_comb begin
    // Default values
    pslverr = 1'b0;
    prdata  = 32'd0;
    if (psel & penable & ~pwrite) begin
      case (paddr)
        ADDR_WDT_CTRL:     prdata = reg_wdt_ctrl;
        ADDR_WDT_TIMEOUT:  prdata = reg_wdt_timeout;
        ADDR_WDT_STATUS:   prdata = reg_wdt_status;
        ADDR_WDT_INT_EN:   prdata = reg_wdt_int_en;
        ADDR_WDT_INT_STAT: prdata = reg_wdt_int_stat;
        default:           pslverr = 1'b1;
      endcase
    end
  end

  // The APB slave is always ready in this design.
  assign pready = 1'b1;

  //-------------------------------------------------------------------------
  // Watchdog Counter Logic (clock gated if enabled)
  //-------------------------------------------------------------------------
  always_ff @(posedge clk_counter or negedge presetn) begin
    if (!presetn) begin
      counter <= 32'd0;
    end else if (reg_wdt_ctrl[CTRL_ENABLE]) begin
      // Check for debug mode pause (if enabled in control register)
      if (reg_wdt_ctrl[CTRL_DEBUG_PAUSE] && debug_mode) begin
        counter <= counter; // Pause counter increment in debug mode
      end
      // Feed event resets the counter if within valid window (or if window mode is disabled)
      else if (feed_event) begin
        counter <= 32'd0;
      end
      // Increment the counter until it reaches the timeout value
      else if (counter < reg_wdt_timeout) begin
        counter <= counter + 1;
      end else begin
        // Once timeout is reached, hold the counter (reset generation is handled below)
        counter <= counter;
      end
    end else begin
      // If watchdog is disabled, keep counter at zero.
      counter <= 32'd0;
    end
  end

  //-------------------------------------------------------------------------
  // Interrupt and Reset Generation Logic (synchronous to pclk)
  //-------------------------------------------------------------------------
  always_ff @(posedge pclk or negedge presetn) begin
    if (!presetn) begin
      reg_wdt_status[0]   <= 1'b0; // Clear timeout status flag
      wdt_reset           <= 1'b0;
      wdt_int             <= 1'b0;
      reg_wdt_int_stat[0] <= 1'b0;
    end else if (reg_wdt_ctrl[CTRL_ENABLE]) begin
      // Generate a pre-timeout interrupt when the counter reaches (timeout - margin)
      if ((counter == (reg_wdt_timeout - INT_MARGIN)) && reg_wdt_int_en[0])
        reg_wdt_int_stat[0] <= 1'b1;
      // Update the external interrupt signal from the interrupt status flag
      wdt_int <= reg_wdt_int_stat[0];

      // If the counter reaches or exceeds the configured timeout, set the status flag and assert reset.
      if (counter >= reg_wdt_timeout) begin
        reg_wdt_status[0] <= 1'b1;
        wdt_reset         <= 1'b1;  // Assert reset (could be a pulse in a real system)
      end else begin
        reg_wdt_status[0] <= 1'b0;
        wdt_reset         <= 1'b0;
      end
    end else begin
      // When WDT is disabled
      reg_wdt_status[0]   <= 1'b0;
      wdt_reset           <= 1'b0;
      wdt_int             <= 1'b0;
      reg_wdt_int_stat[0] <= 1'b0;
    end
  end

endmodule
